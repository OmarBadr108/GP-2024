/*//////////////////////////////////////////////////////////////////////////////////
==================================================================================
 MIXEL GP 2024 LIBRARY
 Copyright (c) 2023 Mixel, Inc.  All Rights Reserved.
 CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF MIXEL and ASU 2024 GP, INC.

 Authors: 
 
 Revision:   

 Version : 1.0

 Create Date: 
 Design Name:  
 Module Name:  

==================================================================================

  STATEMENT OF USE

  This information contains confidential and proprietary information of MIXEL.
  No part of this information may be reproduced, transmitted, transcribed,
  stored in a retrieval system, or translated into any human or computer
  language, in any form or by any means, electronic, mechanical, magnetic,
  optical, chemical, manual, or otherwise, without the prior written permission
  of MIXEL.  This information was prepared for Garduation Project purpose and is for
  use by MIXEL Engineers only.  MIXEL and ASU 2023 GP reserves the right 
  to make changes in the information at any time and without notice.

==================================================================================
//////////////////////////////////////////////////////////////////////////////////*/

module RX (

input                     i_sys_clk,
input                     i_sys_rst,
input                     i_sclgen_scl,
input                     i_sclgen_scl_pos_edge,
input                     i_sclgen_scl_neg_edge,
input                     i_ddrccc_rx_en,
input                     i_sdahnd_rx_sda,
input     [4:0]           i_bitcnt_rx_bit_count,
input     [2:0]           i_ddrccc_rx_mode,
input                     i_crc_value,
input                     i_crc_valid,

output    [7:0]           o_regfcrc_rx_data_out,
output                    o_ddrccc_rx_mode_done,
output                    o_ddrccc_second_pre,
output                    o_ddrccc_error,
output                    o_crc_en                 

);

///////////rx modes///////////

localparam [3:0]  
                     PREAMBLE            = 4'b0000  , 
                     NACK_BIT            = 4'b0001  ,        
                     Deserializing_byte  = 'b0011 ,                   
                     Check_token         = 'b0101 ,
                     Check_Parity_value  = 'b0110 ,
                     Check_CRC_value     = 'b0111 ,
                     Error               = 'b1000 ;










  );
endmodule