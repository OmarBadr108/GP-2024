/*//////////////////////////////////////////////////////////////////////////////////
==================================================================================
 MIXEL GP 2024 LIBRARY
 Copyright (c) 2023 Mixel, Inc.  All Rights Reserved.
 CONFIDENTIAL AND PROPRIETARY SOFTWARE/DATA OF MIXEL and ASU 2024 GP, INC.

 Authors: Fatma Saad Abdallah
 
 Revision:   

 Version : 1.0

 Create Date: 18/2/2024
 Design Name:  HDR_ENGINE
 Module Name:  hdr_engine

==================================================================================

  STATEMENT OF USE

  This information contains confidential and proprietary information of MIXEL.
  No part of this information may be reproduced, transmitted, transcribed,
  stored in a retrieval system, or translated into any human or computer
  language, in any form or by any means, electronic, mechanical, magnetic,
  optical, chemical, manual, or otherwise, without the prior written permission
  of MIXEL.  This information was prepared for Garduation Project purpose and is for
  use by MIXEL Engineers only.  MIXEL and ASU 2023 GP reserves the right 
  to make changes in the information at any time and without notice.

==================================================================================
//////////////////////////////////////////////////////////////////////////////////*/
module hdr_engine (
    input   wire            i_sys_clk                             ,
    input   wire            i_sys_rst_n                           ,
    input   wire            i_i3cengine_hdrengine_en              , 
    input   wire            i_ccc_done                            ,
    input   wire            i_ddr_mode_done                       ,
    input   wire            i_TOC                                 , //term of completion if 0 restart/ 1 exit needed for exit
    input   wire            i_CP                                  , // Cmnd present=1 if CCC 0 for Normal Transcation
    //input   wire  [3:0]     i_TID                                 , //Transaction id for each CCC
    input   wire  [2:0]     i_MODE                                ,
    //to_blocks
    output  reg             o_i3cengine_hdrengine_done            ,
    output  reg             o_ddrmode_en                          ,
    output  reg             o_ccc_en                              ,
    output  reg   [7:0]     o_regf_addr_special
    //config
    //output  reg   [3:0]     o_TID                                 ,
    //output  reg   [7:0]     o_ERR_STATUS                          ,
    //output  reg   [15:0]    o_DATA_LENGTH                         

    );
/////////////parameters////////////
localparam  IDLE          = 2'b00;
localparam  CCC           = 2'b01;
localparam  DDR_MODE      = 2'b10;

reg current_state, next_state;
reg ccc_done;

//--------------------------------- main ------------------------------------------------

always @(posedge i_sys_clk or negedge i_sys_rst_n ) 
  begin: hdr_engine_fsm
    if (!i_sys_rst_n) 
        begin
            o_i3cengine_hdrengine_done      <= 1'b0   ;
            o_hdrmode_en                    <= 1'b0   ;
            o_ccc_en                        <= 1'b0   ;
            o_regf_addr_special             <= 8'd10000 ;
            current_state                   <= IDLE ;
        end

    else if (i_i3cengine_hdrengine_en)
      begin
        current_state <= next_state;
        case (current_state)
          IDLE : begin
              if(i_CP) begin
                  o_ccc_en        <= 1'b1 ;
                  next_state      <= CCC ;
                end
              else 
              begin
                o_ddrmode_en      <= 1'b1 ;
                next_state        <= DDR_MODE ;
              end
          end
          CCC : begin
            if((i_TOC && i_ccc_done)||(i_MODE != 'd6)) begin
                  o_ccc_en    <= 1'b0 ;
                  ccc_done <= 1'b1 ;

                  if(!i_CP) 
                  begin
                    ccc_done <= 1'b0 ;
                    o_regf_addr_special <= 8'd900; //go to special address to get dummy value
                    o_ccc_en   <= 1'b1 ;
                    next_state <= CCC ;
                  end
                  else
                    next_state <= CCC ;

                  if(!i_CP && ccc_done)
                    next_state <= DDR_MODE ;
                  else
                    o_i3cengine_hdrengine_done      <= 1'b1 ;
            end
            else
                  o_i3cengine_hdrengine_done      <= 1'b0 ;
          end
          DDR_MODE : begin
            if ((i_TOC && i_ddr_mode_done)||(i_MODE != 'd6)) begin
              o_ddrmode_en    <= 1'b0 ;
              o_i3cengine_hdrengine_done      <= 1'b1 ;
            end
            else
              begin
                o_ddrmode_en    <= 1'b1 ;
                o_i3cengine_hdrengine_done      <= 1'b0 ;
              end
          end
        endcase
      end

        
end 
endmodule



/*begin
            if (i_i3cengine_hdrengine_en) 
            begin
                if(i_CP) begin
                    o_ccc_en        <= 1'b1 ;
                    if((i_TOC && i_ccc_done)||(i_MODE != 'd6)) begin
                        o_ccc_en    <= 1'b0 ;
                        o_i3cengine_hdrengine_done      <= 1'b1 ;
                      end
                    else
                        o_i3cengine_hdrengine_done      <= 1'b0 ;
                end
                else if (!i_CP) 
                begin
                    o_hdrmode_en        <= 1'b1 ;
                    if((i_TOC && i_hdr_mode_done)||(i_MODE != 'd6)) begin
                        o_hdrmode_en    <= 1'b0 ;
                        o_i3cengine_hdrengine_done      <= 1'b1 ;
                      end
                    else
                        o_i3cengine_hdrengine_done      <= 1'b0 ;
                end
                else begin
                  o_i3cengine_hdrengine_done      <= 1'b0 ;
                  o_ccc_en                        <= 1'b0  ;
                  o_hdrmode_en                    <= 1'b0  ; 
                end
            end
            else
                begin
                    o_i3cengine_hdrengine_done      <= 1'b0  ;
                    o_ccc_en                        <= 1'b0  ;
                    o_hdrmode_en                    <= 1'b0  ;

                end

            
        end*/
